moduele();
endmodule;
